`ifndef _bp_
`define _bp_

class Basepacket;
	randc logic[3:0]i;
	logic en;
	logic [15:0]y;
endclass : Basepacket

`endif