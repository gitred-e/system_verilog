`ifndef _bp_
`define _bp_

class Basepacket;
	bit rst;
	bit [3:0]q;
endclass : Basepacket

`endif