module dec_design(dec_intf.dec_dut intf);

	always @(*) begin
		if(intf.en) begin
			case(intf.i)
				'd0:begin
					intf.y[0]='b1;
					intf.y[15:1]='b0;
				end
				'd1:begin
					intf.y[1]='b1;
					intf.y[0]='b0;
					intf.y[15:2]='b0;
				end
				'd2:begin
					intf.y[2]='b1;
					intf.y[1:0]='b0;
					intf.y[15:3]='b0;
				end
				'd3:begin
					intf.y[3]='b1;
					intf.y[2:0]='b0;
					intf.y[15:4]='b0;
				end
				'd4:begin
					intf.y[4]='b1;
					intf.y[3:0]='b0;
					intf.y[15:5]='b0;
				end
				'd5:begin
					intf.y[5]='b1;
					intf.y[4:0]='b0;
					intf.y[15:6]='b0;
				end
				'd6:begin
					intf.y[6]='b1;
					intf.y[5:0]='b0;
					intf.y[15:7]='b0;
				end
				'd7:begin
					intf.y[7]='b1;
					intf.y[6:0]='b0;
					intf.y[15:8]='b0;
				end
				'd8:begin
					intf.y[8]='b1;
					intf.y[7:0]='b0;
					intf.y[15:9]='b0;
				end
				'd9:begin
					intf.y[9]='b1;
					intf.y[8:0]='b0;
					intf.y[15:10]='b0;
				end
				'd10:begin
					intf.y[10]='b1;
					intf.y[9:0]='b0;
					intf.y[15:11]='b0;
				end
				'd11:begin
					intf.y[11]='b1;
					intf.y[10:0]='b0;
					intf.y[15:12]='b0;
				end
				'd12:begin
					intf.y[12]='b1;
					intf.y[11:0]='b0;
					intf.y[15:13]='b0;
				end
				'd13:begin
					intf.y[13]='b1;
					intf.y[12:0]='b0;
					intf.y[15:14]='b0;
				end
				'd14:begin
					intf.y[14]='d1;
					intf.y[13:0]='d0;
					intf.y[15]='d0;
				end
				'd15:begin
					intf.y[15]='b1;
					intf.y[14:0]='b0;
				end
				default:intf.y='bx;
			endcase // intf.i
		end
		else
			intf.y='b0;
	end
endmodule : dec_design